library verilog;
use verilog.vl_types.all;
entity frame_gen_tb is
end frame_gen_tb;
