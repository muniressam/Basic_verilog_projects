library verilog;
use verilog.vl_types.all;
entity baudGen_tb is
end baudGen_tb;
