library verilog;
use verilog.vl_types.all;
entity piso_tb is
end piso_tb;
